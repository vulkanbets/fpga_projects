`timescale 1ns / 1ns

module hello
(
    input A,
    output wire B
);

    assign B = A;

endmodule
