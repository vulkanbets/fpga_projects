`timescale 1ns / 1ns

module hello
(
    input A,
    output B
);

    assign B = A;

endmodule
